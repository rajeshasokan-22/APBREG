`ifndef DUT_WRAPPER_SV
`define DUT_WRAPPER_SV

`include "uvm_macros.svh"
import uvm_pkg::*;

module dut_wrapper();
    
endmodule

`endif

